package PacketTest;
import NocPacket::*;
import Packet::*;


module mkPacketTest();       
   rule hello;
      $finish;                   
   endrule
endmodule
endpackage